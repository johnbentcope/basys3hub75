module HUB75Driver(output [7:0] JB, JC, input clk);

  reg A0, A1, A2, A3, A4, BL, CK, LA, R0, G0, B0, R1, G1, B1, X0, X1;

  assign A0 = rowCounterLow[0];
  assign A1 = rowCounterLow[1];
  assign A2 = rowCounterLow[2];
  assign A3 = 0;
  assign A4 = 0;

  assign JB = {R0, G0, B0, X0, R1, G1, B1, X1};
  assign JC = {A0, A1, A2, A3, BL, LA, CK, A4};

  reg [32:0] clockCounter;
  reg [2:0] rowCounterLow <= 0;
  reg [3:0] rowCounterHigh;
  assign rowCounterHigh = {{1{1}}, rowCounterLow}; // Will always move lock-step with the other
  reg [4:0] columnCounter;

  wire pixelClock;
  
  // NOT PERMANENT DATA. TEST DATA WHILE TIMING BUILT
  reg [31:0]red[15:0];
  reg [31:0]grn[15:0];
  reg [31:0]blu[15:0];
  red[0] = 32'b01010101_01010101_01010101_01010101;
  red[1] = 32'b01010101_01010101_01010101_01010101;
  red[2] = 32'b01010101_01010101_01010101_01010101;
  red[3] = 32'b01010101_01010101_01010101_01010101;
  red[4] = 32'b00110011_00110011_00110011_00110011;
  red[5] = 32'b00110011_00110011_00110011_00110011;
  red[6] = 32'b00110011_00110011_00110011_00110011;
  red[7] = 32'b00110011_00110011_00110011_00110011;
  red[8] = 32'b00001111_00001111_00001111_00001111;
  red[9] = 32'b00001111_00001111_00001111_00001111;
  red[10] = 32'b00001111_00001111_00001111_00001111;
  red[11] = 32'b00001111_00001111_00001111_00001111;
  red[12] = 32'b00000000_11111111_00000000_11111111;
  red[13] = 32'b00000000_11111111_00000000_11111111;
  red[14] = 32'b00000000_11111111_00000000_11111111;
  red[15] = 32'b00000000_11111111_00000000_11111111;
  grn[0] = 32'b00110011_00110011_00110011_00110011;
  grn[1] = 32'b00110011_00110011_00110011_00110011;
  grn[2] = 32'b00110011_00110011_00110011_00110011;
  grn[3] = 32'b00110011_00110011_00110011_00110011;
  grn[4] = 32'b00001111_00001111_00001111_00001111;
  grn[5] = 32'b00001111_00001111_00001111_00001111;
  grn[6] = 32'b00001111_00001111_00001111_00001111;
  grn[7] = 32'b00001111_00001111_00001111_00001111;
  grn[8] = 32'b00000000_11111111_00000000_11111111;
  grn[9] = 32'b00000000_11111111_00000000_11111111;
  grn[10] = 32'b00000000_11111111_00000000_11111111;
  grn[11] = 32'b00000000_11111111_00000000_11111111;
  grn[12] = 32'b01010101_01010101_01010101_01010101;
  grn[13] = 32'b01010101_01010101_01010101_01010101;
  grn[14] = 32'b01010101_01010101_01010101_01010101;
  grn[15] = 32'b01010101_01010101_01010101_01010101;
  blu[0] = 32'b00001111_00001111_00001111_00001111;
  blu[1] = 32'b00001111_00001111_00001111_00001111;
  blu[2] = 32'b00001111_00001111_00001111_00001111;
  blu[3] = 32'b00001111_00001111_00001111_00001111;
  blu[4] = 32'b00000000_11111111_00000000_11111111;
  blu[5] = 32'b00000000_11111111_00000000_11111111;
  blu[6] = 32'b00000000_11111111_00000000_11111111;
  blu[7] = 32'b00000000_11111111_00000000_11111111;
  blu[8] = 32'b01010101_01010101_01010101_01010101;
  blu[9] = 32'b01010101_01010101_01010101_01010101;
  blu[10] = 32'b01010101_01010101_01010101_01010101;
  blu[11] = 32'b01010101_01010101_01010101_01010101;
  blu[12] = 32'b00110011_00110011_00110011_00110011;
  blu[13] = 32'b00110011_00110011_00110011_00110011;
  blu[14] = 32'b00110011_00110011_00110011_00110011;
  blu[15] = 32'b00110011_00110011_00110011_00110011;
  
w
  initial
  begin
    BL <= 0;
    LA <= 0;
    CK <= 0;

    R0 <= 0;
    R1 <= 1;
    G0 <= 0;
    G1 <= 1;
    B0 <= 0;
    B1 <= 1;
    X0 <= 0;
    X1 <= 0;
    clockCounter <= 0;
  end

  // States
  // Shifting out data loop
  // Blank display
  // Latch data
  // Unblank display and increment address

  reg [1:0] CS, NS;

  always @(posedge clk)
  begin
    clockCounter <= clockCounter + 1;
    case(CS)
      0: NS <= (clockCounter < 32) CS : NS;
    endcase
  end

endmodule